--
-- TCPA VHDL code generator
--
-- File: wppa_top.vhd
-- Date: 30.05.2017
-- Time: 14:38:13
--

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

library wppa_instance_v1_01_a;
use wppa_instance_v1_01_a.ALL;
use wppa_instance_v1_01_a.WPPE_LIB.ALL;
use wppa_instance_v1_01_a.DEFAULT_LIB.ALL;
use wppa_instance_v1_01_a.ARRAY_LIB.ALL;
use wppa_instance_v1_01_a.TYPE_LIB.ALL;
use wppa_instance_v1_01_a.INVASIC_LIB.all;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


-- Entity port declaration with input and output signals of
-- WPPA model and implicitly clock and asynchronous reset

ENTITY WPPA_TOP IS

	GENERIC(
					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%

					 -- cadence translate_off 
					 INSTANCE_NAME                  :string := "TOP_LEVEL_MODULE";
					 -- cadence translate_on 
					 wppa_generics  :t_wppa_generics := DEFAULT_WPPA_GENERICS 
		);

	PORT(
					--/////////////////////////////////////////////////--

                clk, rst                     : in  std_logic;

                -- Bus 
                wppa_bus_input_interface     : in  t_wppa_bus_input_interface;
                wppa_bus_output_interface    : out t_wppa_bus_output_interface;
                -- Data 
                wppa_data_input              : in  t_wppa_data_input_interface;
                wppa_data_output             : out t_wppa_data_output_interface;
                -- Control 
                wppa_ctrl_input              : in  t_wppa_ctrl_input_interface;
                wppa_ctrl_output             : out t_wppa_ctrl_output_interface;
                wppa_memory_input_interface  : in  t_wppa_memory_input_interface;
                wppa_memory_output_interface : out t_wppa_memory_output_interface;
                fault_injection              : in  t_fault_injection_module;
                error_status                 : out t_error_status;
                tcpa_config_done             : out std_logic;
                tcpa_config_done_vector      : out std_logic_vector(31 downto 0);
                ctrl_programmable_depth      : in  t_ctrl_programmable_depth;
                en_programmable_fd_depth     : in  t_en_programmable_fd_depth;
                programmable_fd_depth        : in  t_programmable_fd_depth;
                enable_tcpa                  : in  std_logic;
                pc_debug_out                 : out t_pc_debug_outs;
                icp_program_interface        : in  t_prog_intfc;
                invasion_input               : in  t_inv_sig;
                invasion_output              : out t_inv_sig;
                parasitary_invasion_input    : in  t_inv_sig;
                parasitary_invasion_output   : out t_inv_sig

		);

END WPPA_TOP;

ARCHITECTURE Behavioral OF WPPA_TOP IS
signal fault_injection_sig : t_fault_injection_module;	

COMPONENT WPPA is

	GENERIC(
					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%

					 -- cadence translate_off 
					 INSTANCE_NAME         :string;
					 WPPA_SIZE             :string;
					 -- cadence translate_on
					 wppa_generics :t_wppa_generics := DEFAULT_WPPA_GENERICS;

					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
					-- GENERICS FOR THE WP PROCESSORS AND THEIR INTERCONNECT WRAPPERS
					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
					------------------------------------------
					ADJ_MATRIX_ARRAY_ALL:t_adj_matrix_array_all(1 to  4, 1 to 4);
					------------------------------------------
					WPPE_GENERICS:t_wppe_generics_array(1 to 4, 1 to 4) 
					------------------------------------------
		);

	PORT(
					--/////////////////////////////////////////////////--

		clk_in, rst                     : in  std_logic;

		-- Bus 
		wppa_bus_input_interface     : in  t_wppa_bus_input_interface;
		wppa_bus_output_interface    : out t_wppa_bus_output_interface;
		-- Data 
		wppa_data_input              : in  t_wppa_data_input_interface;
		wppa_data_output             : out t_wppa_data_output_interface;
		-- Control 
		wppa_ctrl_input              : in  t_wppa_ctrl_input_interface;
		wppa_ctrl_output             : out t_wppa_ctrl_output_interface;
		wppa_memory_input_interface  : in  t_wppa_memory_input_interface;
		wppa_memory_output_interface : out t_wppa_memory_output_interface;
		fault_injection              : in  t_fault_injection_module;
		error_status                 : out t_error_status; 
		tcpa_config_done             : out std_logic;
		tcpa_config_done_vector      : out std_logic_vector(31 downto 0);
		ctrl_programmable_depth      : in  t_ctrl_programmable_depth;
		en_programmable_fd_depth     : in  t_en_programmable_fd_depth;
		programmable_fd_depth        : in  t_programmable_fd_depth;
		enable_tcpa                  : in  std_logic;
		pc_debug_out                 : out t_pc_debug_outs;		
		icp_program_interface        : in  t_prog_intfc;
		invasion_input               : in  t_inv_sig;
		invasion_output              : out t_inv_sig;
		parasitary_invasion_input    : in  t_inv_sig;
		parasitary_invasion_output   : out t_inv_sig

		);

END COMPONENT;

BEGIN


internal_wppa :WPPA

	generic map(
					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%

					-- cadence translate_off
					INSTANCE_NAME => "wppa_top",
					WPPA_SIZE     => "4x4",
					-- cadence translate_on
					wppa_generics => wppa_generics,

					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
					-- GENERICS FOR THE WP PROCESSORS AND THEIR INTERCONNECT WRAPPERS
					--%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
					------------------------------------------
					ADJ_MATRIX_ARRAY_ALL  	   =>	(
					--==============================================================
					--==============================================================
------------------------
(  --     0. WPPA ROW
------------------------
-- P[0,0] ADJ_MATRIX
( "0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[0,1] ADJ_MATRIX
( "0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000001111100000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[0,2] ADJ_MATRIX
( "0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000001111100000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[0,3] ADJ_MATRIX
( "0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000001111100000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
)
),--     END0. WPPA ROW
------------------------
(  --     1. WPPA ROW
------------------------
-- P[1,0] ADJ_MATRIX
( "0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[1,1] ADJ_MATRIX
( "0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000001111100000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[1,2] ADJ_MATRIX
( "0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000001111100000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[1,3] ADJ_MATRIX
( "0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000001111100000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
)
),--     END1. WPPA ROW
------------------------
(  --     2. WPPA ROW
------------------------
-- P[2,0] ADJ_MATRIX
( "0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[2,1] ADJ_MATRIX
( "0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000001111100000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[2,2] ADJ_MATRIX
( "0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000001111100000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[2,3] ADJ_MATRIX
( "0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000001111100000000000000",
"0000000000000000000000000000010",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"1111001111101111001111000000000",
"0000000000100000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
)
),--     END2. WPPA ROW
------------------------
(  --     3. WPPA ROW
------------------------
-- P[3,0] ADJ_MATRIX
( "0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"0000000000000000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[3,1] ADJ_MATRIX
( "0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"0000000000000000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[3,2] ADJ_MATRIX
( "0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"0000000000000000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
),
-- P[3,3] ADJ_MATRIX
( "0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000001111100",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000001111000",
"0000000000000000000000000000000",
"0000000000000000000000000000010",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"1111001111001111001111000000000",
"0000000000000000000000000000000",
"0000010000010000010000010000000",
"0000000000000000000000000000000"
)
)--     END3. WPPA ROW
												--==============================================================
													--==============================================================	
													),

					------------------------------------------
					WPPE_GENERICS 	  			=>	(
					------------------------------------------
					 (  -- BEGIN WPPA 0 ROW
					     --##############################################################################
					  ( -- BEGIN WPPE[0,0] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[0,0] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[0,1] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[0,1] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[0,2] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[0,2] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[0,3] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  )  -- END WPPE[0,3] GENERICS RECORD
					     --##############################################################################

					 ), -- END WPPA 0 ROW
					 (  -- BEGIN WPPA 1 ROW
					     --##############################################################################
					  ( -- BEGIN WPPE[1,0] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[1,0] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[1,1] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[1,1] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[1,2] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[1,2] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[1,3] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  )  -- END WPPE[1,3] GENERICS RECORD
					     --##############################################################################

					 ), -- END WPPA 1 ROW
					 (  -- BEGIN WPPA 2 ROW
					     --##############################################################################
					  ( -- BEGIN WPPE[2,0] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[2,0] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[2,1] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[2,1] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[2,2] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[2,2] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[2,3] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  )  -- END WPPE[2,3] GENERICS RECORD
					     --##############################################################################

					 ), -- END WPPA 2 ROW
					 (  -- BEGIN WPPA 3 ROW
					     --##############################################################################
					  ( -- BEGIN WPPE[3,0] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[3,0] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[3,1] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[3,1] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[3,2] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  ), -- END WPPE[3,2] GENERICS RECORD
					     --##############################################################################

					     --##############################################################################
					  ( -- BEGIN WPPE[3,3] GENERICS RECORD
					     --##############################################################################

										CUR_DEFAULT_CONFIG_REG_WIDTH,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF BRANCH FLAGS
										--*******************************************************************************--

										2,

										--*****************************************************************************************--
										-- GENERICS FOR THE NUMBER OF CONTROL REGISTERS, CONTROL INPUTS and CONTROL OUTPUTS
										--*****************************************************************************************--

										1,
										2,
										2,

										--*******************************************************************************--
										-- GENERICS FOR THE CONTROL REGISTER WIDTH --
										--*******************************************************************************--

										1,

										--*******************************************************************************--
										-- GENERICS FOR THE CTRL REGISTERS ADDRESS WIDTH
										--*******************************************************************************--

										5, -- RegField Width

										--*******************************************************************************--
										-- GENERICS FOR CONFIGURATION MEMORY
										--*******************************************************************************--

										CUR_DEFAULT_SOURCE_ADDR_WIDTH,
										CUR_DEFAULT_SOURCE_DATA_WIDTH,

										--*******************************************************************************--
										-- Turning the ASSERT ... messages on for simulation and off for synthesis
										--*******************************************************************************--

										--					CUR_DEFAULT_SIMULATION,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT INSTRUCTION WIDTH
										--*******************************************************************************--

										18,

										--*******************************************************************************--
										-- GENERICS FOR THE CURRENT BRANCH INSTRUCTION WIDTH
										--*******************************************************************************--

										49,

										--*******************************************************************************--
										-- GENERICS FOR THE INSTRUCTION MEMORY SIZE
										--*******************************************************************************--

										96,

										--*******************************************************************************--
										-- GENERICS FOR THE ADDRESS AND DATA WIDTHS
										--*******************************************************************************--

										7, -- InstrMem Addr Width 
										5, -- RegField Width
										32, -- Data Path Width

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF SPECIFIC FUNCTIONAL UNITS
										--*******************************************************************************--

										2, -- Adders Number 
										1,  -- Mult Number 
										0,   -- Div Number 
										1, -- LogicFU Number 
										1, -- ShiftFU Number 
										6,   -- DPU Number 
										2,   -- CPU Number 


										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF INPUT AND OUTPUT REGISTERS 
										--*******************************************************************************--

										5, -- NumOf Output Regs 
										5,  -- NumOf Input Regs 

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER OF THE GENERAL PURPOSE REGISTERS
										--*******************************************************************************--

										16,

										--*******************************************************************************--
										-- GENERICS FOR THE NUMBER AND SIZE OF additional FIFOs --
										--*******************************************************************************--

										3, -- Number FB FIFOs 
										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "111", -- Type FB FIFOs
										(16, 16, 16), -- Size FB FIFOs
										(4, 4, 4), -- Addr width FB FIFOs

										-- When LUT_RAM_TYPE = '1' => LUT_RAM, else BLOCK_RAM
										 "11111", -- TYPE Input FIFOs
										(1, 1, 1, 1, 1), -- Size Input FIFOs
										(1, 1, 1, 1, 1), -- Addr Width Input FIFOs 

										--*******************************************************************************--
										-- GENERICS FOR THE WIDH OF ALL REGISTERS
										--*******************************************************************************--

										32

					     --##############################################################################
					  )  -- END WPPE[3,3] GENERICS RECORD
					     --##############################################################################

					 )  -- END WPPA 3 ROW
					) -- END WPPA ARRAY
	)   -- END GENERIC MAP
	PORT MAP(

			--/////////////////////////////////////////////////--

                        clk_in                       => clk,
                        rst                          => rst,

                        -- Bus
                        wppa_bus_input_interface     => wppa_bus_input_interface,
                        wppa_bus_output_interface    => wppa_bus_output_interface,
                        -- Data
                        wppa_data_input              => wppa_data_input,
                        wppa_data_output             => wppa_data_output,
                        -- Control
                        wppa_ctrl_input              => wppa_ctrl_input,
                        wppa_ctrl_output             => wppa_ctrl_output,
                        -- Memory
                        wppa_memory_input_interface  => wppa_memory_input_interface,
                        wppa_memory_output_interface => wppa_memory_output_interface,
                        tcpa_config_done             => tcpa_config_done,
                        fault_injection              => fault_injection_sig,	
                        error_status                  => error_status,
                        tcpa_config_done_vector      => tcpa_config_done_vector,
                        ctrl_programmable_depth      => ctrl_programmable_depth,
                        en_programmable_fd_depth     => en_programmable_fd_depth,
                        programmable_fd_depth        => programmable_fd_depth,
                        enable_tcpa                  => enable_tcpa,
                        pc_debug_out                 => pc_debug_out,
                        icp_program_interface        => icp_program_interface,
                        invasion_input               => invasion_input,
                        invasion_output              => invasion_output,
                        parasitary_invasion_input    => parasitary_invasion_input,
                        parasitary_invasion_output   => parasitary_invasion_output
	);

	sync : process(clk)
	begin
		if rising_edge(clk) then

				fault_injection_sig.mask   <= fault_injection.mask;
				fault_injection_sig.fu_sel <= fault_injection.fu_sel;
				fault_injection_sig.pe_sel <= fault_injection.pe_sel;

		end if;
	end process;


END Behavioral;

