---------------------------------------------------------------------------------------------------------------------------------
-- (C) Copyright 2013 Chair for Hardware/Software Co-Design, Department of Computer Science 12,
-- University of Erlangen-Nuremberg (FAU). All Rights Reserved
--------------------------------------------------------------------------------------------------------------------------------
-- Module Name:  
-- Project Name:  
--
-- Engineer:     
-- Create Date:   
-- Description:  
--
--------------------------------------------------------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:    14:15:08 01/04/06
-- Design Name:    
-- Module Name:    config_memory - Behavioral
-- Project Name:   
-- Target Device:  
-- Tool versions:  
-- Description:
--
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
--------------------------------------------------------------------------------
library IEEE;
library wppa_instance_v1_01_a;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- pragma translate_off
-- cadence translate_on
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use std.textio.all;
use IEEE.std_logic_textio.all;
-- pragma translate_on

library wppa_instance_v1_01_a;
use wppa_instance_v1_01_a.ALL;

use wppa_instance_v1_01_a.WPPE_LIB.all;
use wppa_instance_v1_01_a.DEFAULT_LIB.all;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity config_memory is
	generic(

		-- cadence translate_off                
		INSTANCE_NAME : string   := "";

		-- cadence translate_on                         
		MEM_SIZE      : positive := CUR_DEFAULT_SOURCE_MEM_SIZE;
		DATA_WIDTH    : positive := CUR_DEFAULT_SOURCE_DATA_WIDTH;
		ADDR_WIDTH    : positive := CUR_DEFAULT_SOURCE_ADDR_WIDTH
	);

	port(
		clk       : in  std_logic;
		rst       : in  std_logic;
		cfg_reset : in  std_logic;
		we        : in  std_logic;
		d_in      : in  std_logic_vector(DATA_WIDTH - 1 downto 0);
		addr      : in  std_logic_vector(ADDR_WIDTH - 1 downto 0);
		d_out     : out std_logic_vector(DATA_WIDTH - 1 downto 0)
	);

end config_memory;

architecture Behavioral of config_memory is
	type t_ram is array (0 to MEM_SIZE - 1) of std_logic_vector(DATA_WIDTH - 1 downto 0);

	signal ram : t_ram := (
		"10000000100101111010000101111001", -- 0x0(0)  Domain_0, Type: VLIW, Vert.Mask:2 "10" Horiz.Mask:2 "10",  *** PE[0,0] *** d0 FIR VLIW
		"11111111111111111111111100010111",
		"11111111111111111111111111111111", -- 0x2(2)  0. VLIW 
		"00101100000000001111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x5(5)  1. VLIW 
		"00101010000000001111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x8(8)  2. VLIW 
		"00101010000000011111111111111111",
		"11111111111000111000011100110010",
		"00100000100000010100010000000000", -- 0xB(11)  3. VLIW 
		"11111111111111111111111111111111",
		"11111111111000000000000000110011",
		"11111111111111111111111111111111", -- 0xE(14)  4. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x11(17)  5. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x14(20)  6. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x17(23)  7. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x1A(26)  8. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x1D(29)  9. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x20(32)  10. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x23(35)  11. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x26(38)  12. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x29(41)  13. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x2C(44)  14. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		--________________________________
		--==  Domain0 Header Parsing: [ Type: 1 (VLIW), lastFlag: 0, Next: 47, Vertical Mask: "10", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 2, VLIW end: 47, ICN begin: 511, ICN end: 511 ]
		--================================
		--
		"00001100010101111001001011110001", -- 0x2F(47)  Domain_1, Type: VLIW, Vert.Mask:1 "01" Horiz.Mask:2 "10",  *** PE[0,1] *** d1 FIR VLIW
		"11111111111111111111111100101111",
		"00100000100000010000001011000000", -- 0x31(49)  0. VLIW 
		"11111111111111111000010000100010",
		"11111111111000000000000000000000",
		"11111111111111111111111111111111", -- 0x34(52)  1. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x37(55)  2. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x3A(58)  3. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x3D(61)  4. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x40(64)  5. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x43(67)  6. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x46(70)  7. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x49(73)  8. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x4C(76)  9. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x4F(79)  10. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x52(82)  11. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x55(85)  12. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x58(88)  13. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x5B(91)  14. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		--________________________________
		--==  Domain1 Header Parsing: [ Type: 1 (VLIW), lastFlag: 0, Next: 94, Vertical Mask: "01", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 49, VLIW end: 94, ICN begin: 511, ICN end: 511 ]
		--================================
		--
		"10011000000101110110010001101001", -- 0x5E(94)  Domain_2, Type: VLIW, Vert.Mask:2 "10" Horiz.Mask:1 "01",  *** PE[1,0] *** d2 FIR
		"11111111111111111111111101000110",
		"00100000001000010000010010100000", -- 0x60(96)  0. VLIW 
		"11111111111111111000001010000000",
		"11111111111000000000000000000000",
		"11111111111111111111111111111111", -- 0x63(99)  1. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x66(102)  2. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x69(105)  3. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x6C(108)  4. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x6F(111)  5. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x72(114)  6. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x75(117)  7. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x78(120)  8. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x7B(123)  9. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x7E(126)  10. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x81(129)  11. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x84(132)  12. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x87(135)  13. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x8A(138)  14. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		--________________________________
		--==  Domain2 Header Parsing: [ Type: 1 (VLIW), lastFlag: 0, Next: 141, Vertical Mask: "10", Horizontal Mask: "01",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 96, VLIW end: 141, ICN begin: 511, ICN end: 511 ]
		--================================
		--
		"00100011110101110101010111100001", -- 0x8D(141)  Domain_3, Type: VLIW, Vert.Mask:1 "01" Horiz.Mask:1 "01",  *** PE[1,1] *** d3 FIR
		"11111111111111111111111101011110",
		"00100000100000010000010010100000", -- 0x8F(143)  0. VLIW 
		"11111111111111111111111111111111",
		"11111111111000000000000000000000",
		"11111111111111111111111111111111", -- 0x92(146)  1. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x95(149)  2. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x98(152)  3. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x9B(155)  4. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x9E(158)  5. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xA1(161)  6. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xA4(164)  7. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xA7(167)  8. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xAA(170)  9. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xAD(173)  10. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xB0(176)  11. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xB3(179)  12. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xB6(182)  13. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xB9(185)  14. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		--________________________________
		--==  Domain3 Header Parsing: [ Type: 1 (VLIW), lastFlag: 0, Next: 188, Vertical Mask: "01", Horizontal Mask: "01",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 143, VLIW end: 188, ICN begin: 511, ICN end: 511 ]
		--================================
		--
		"11111111110101111010010111111010", -- 0xBC(188)  Domain_4, Type: ICN, Vert.Mask:2 "10" Horiz.Mask:2 "10",  *** PE[0,0] *** d4 FIR ICN
		"11111101011111101011111011111111",
		"11111111111111111111000000111111",
		--________________________________
		--==  Domain4 Header Parsing: [ Type: 2 (ICN), lastFlag: 0, Next: 191, Vertical Mask: "10", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 511, VLIW end: 511, ICN begin: 190, ICN end: 191 ]
		--================================
		--
		"11111111110101111001011000010110", -- 0xBF(191)  Domain_5, Type: ICN, LAST, Vert.Mask:1 "01" Horiz.Mask:2 "10",  *** PE[0,1] *** d5 FIR ICN
		"11111101100001001100000111111111",
		"11111111111111111111111111000001",
		--________________________________
		--==  Domain5 Header Parsing: [ Type: 2 (ICN), lastFlag: 1, Next: 194, Vertical Mask: "01", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 511, VLIW end: 511, ICN begin: 193, ICN end: 194 ]
		--================================
		--
		"10110001000101111010011110001001", -- 0xC2(194)  Domain_6, Type: VLIW, Vert.Mask:2 "10" Horiz.Mask:2 "10",  *** PE[0,0] *** d0 EDGE
		"11111111111111111111111101111000",
		"11111111111111111111111111111111", -- 0xC4(196)  0. VLIW 
		"00101100000000011111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xC7(199)  1. VLIW 
		"00101010000000001111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xCA(202)  2. VLIW 
		"00101010000000011111111111111111",
		"11111111111000111000011100110010",
		"00100000100111110000010000000010", -- 0xCD(205)  3. VLIW 
		"00101000000000011111111111111111",
		"11111111111111000000000000000000",
		"00100000100111100100001000000000", -- 0xD0(208)  4. VLIW 
		"00101000000000001111111111111111",
		"11111111111111000000000000000000",
		"00100000100111110000001000000010", -- 0xD3(211)  5. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111110000001000000010", -- 0xD6(214)  6. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xD9(217)  7. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"00100000100000011111111111111111", -- 0xDC(220)  8. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"00100000100000100000001000000010", -- 0xDF(223)  9. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"00100000100000010000001000000010", -- 0xE2(226)  10. VLIW 
		"11111111111111111111111111111111",
		"11111111111000000000000000110011",
		"11111111111111111111111111111111", -- 0xE5(229)  11. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xE8(232)  12. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xEB(235)  13. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xEE(238)  14. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		--________________________________
		--==  Domain6 Header Parsing: [ Type: 1 (VLIW), lastFlag: 0, Next: 241, Vertical Mask: "10", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 196, VLIW end: 241, ICN begin: 511, ICN end: 511 ]
		--================================
		--
		"00111100110101111001100100000001", -- 0xF1(241)  Domain_7, Type: VLIW, Vert.Mask:1 "01" Horiz.Mask:2 "10",  *** PE[0,1] *** d1 EDGE
		"11111111111111111111111110010000",
		"11111111111111111111111111111111", -- 0xF3(243)  0. VLIW 
		"11111111111111111111111111111111",
		"11111111111000111000011100010000",
		"11111111111111110100000010100000", -- 0xF6(246)  1. VLIW 
		"11111111111111111111111111111111",
		"11111111111000000010000000100011",
		"00100000000111111111111111111111", -- 0xF9(249)  2. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0xFC(252)  3. VLIW 
		"11111111111111111111111111111111",
		"11111111111000111000100001000011",
		"11111111111111110000000000001100", -- 0xFF(255)  4. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x102(258)  5. VLIW 
		"11111111111111111000010000000010",
		"11111111111000000000000000000000",
		"11111111111111111111111111111111", -- 0x105(261)  6. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x108(264)  7. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x10B(267)  8. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x10E(270)  9. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x111(273)  10. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x114(276)  11. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x117(279)  12. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x11A(282)  13. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x11D(285)  14. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		--________________________________
		--==  Domain7 Header Parsing: [ Type: 1 (VLIW), lastFlag: 0, Next: 288, Vertical Mask: "01", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 243, VLIW end: 288, ICN begin: 511, ICN end: 511 ]
		--================================
		--
		"11001000100101110110101001111001", -- 0x120(288)  Domain_8, Type: VLIW, Vert.Mask:2 "10" Horiz.Mask:1 "01",  *** PE[1,0] *** d2 EDGE
		"11111111111111111111111110100111",
		"11111111111111111111111111111111", -- 0x122(290)  0. VLIW 
		"11111111111111111111111111111111",
		"11111111111000111000011100010000",
		"00100000100111110000010000000010", -- 0x125(293)  1. VLIW 
		"00101000000000011111111111111111",
		"11111111111111000000000000000000",
		"11111111111111110100001000000000", -- 0x128(296)  2. VLIW 
		"00101000000000001111111111111111",
		"11111111111111000000000000000000",
		"00100000100000011111111111111111", -- 0x12B(299)  3. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"00100000100111100000001000000010", -- 0x12E(302)  4. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"00100000100000100000001000000010", -- 0x131(305)  5. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"00100000100111110000001000000010", -- 0x134(308)  6. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111110000001000000010", -- 0x137(311)  7. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"00100000100000011111111111111111", -- 0x13A(314)  8. VLIW 
		"11111111111111111111111111111111",
		"11111111111000000000000000010001",
		"11111111111111111111111111111111", -- 0x13D(317)  9. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x140(320)  10. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x143(323)  11. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x146(326)  12. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x149(329)  13. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x14C(332)  14. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		--________________________________
		--==  Domain8 Header Parsing: [ Type: 1 (VLIW), lastFlag: 0, Next: 335, Vertical Mask: "10", Horizontal Mask: "01",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 290, VLIW end: 335, ICN begin: 511, ICN end: 511 ]
		--================================
		--
		"01010100010101110101101111110001", -- 0x14F(335)  Domain_9, Type: VLIW, Vert.Mask:1 "01" Horiz.Mask:1 "01",  *** PE[1,1] *** d3 EDGE VLIW
		"11111111111111111111111110111111",
		"11111111111111111111111111111111", -- 0x151(337)  0. VLIW 
		"00101000000000101111111111111111",
		"11111111111000111000011100010000",
		"11111111111111110100000010100000", -- 0x154(340)  1. VLIW 
		"11111111111111111111111111111111",
		"11111111111000000010000000100011",
		"00100000000111111111111111111111", -- 0x157(343)  2. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111110100010000000000", -- 0x15A(346)  3. VLIW 
		"00101000000000011111111111111111",
		"11111111111000000000000000000000",
		"11111111111111111111111111111111", -- 0x15D(349)  4. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x160(352)  5. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x163(355)  6. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x166(358)  7. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x169(361)  8. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x16C(364)  9. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x16F(367)  10. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x172(370)  11. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x175(373)  12. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x178(376)  13. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x17B(379)  14. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		--________________________________
		--==  Domain9 Header Parsing: [ Type: 1 (VLIW), lastFlag: 0, Next: 382, Vertical Mask: "01", Horizontal Mask: "01",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 337, VLIW end: 382, ICN begin: 511, ICN end: 511 ]
		--================================
		--
		"11111111110101111010110000001010", -- 0x17E(382)  Domain_10, Type: ICN, Vert.Mask:2 "10" Horiz.Mask:2 "10",  *** PE[0,0] *** d4 EDGE ICN
		"11111111000000111000000011111111",
		"11111111111111111111000001111111",
		--________________________________
		--==  Domain10 Header Parsing: [ Type: 2 (ICN), lastFlag: 0, Next: 385, Vertical Mask: "10", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 511, VLIW end: 511, ICN begin: 384, ICN end: 385 ]
		--================================
		--
		"11111111110101111001110000100110", -- 0x181(385)  Domain_11, Type: ICN, LAST, Vert.Mask:1 "01" Horiz.Mask:2 "10",  *** PE[0,1] *** d5 EDGE ICN
		"11111111000010011000001111111111",
		"11111111111111111111111111000001",
		--________________________________
		--==  Domain11 Header Parsing: [ Type: 2 (ICN), lastFlag: 1, Next: 388, Vertical Mask: "01", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 511, VLIW end: 511, ICN begin: 387, ICN end: 388 ]
		--================================
		--
		"11100001100101111010110110011001", -- 0x184(388)  Domain_12, Type: VLIW, Vert.Mask:2 "10" Horiz.Mask:2 "10",  *** PE[0,0] *** d0 INVERT VLIW
		"11111111111111111111111111011001",
		"11111111111111111111111111111111", -- 0x186(390)  0. VLIW 
		"00101100000000001111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x189(393)  1. VLIW 
		"00101010000000001111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x18C(396)  2. VLIW 
		"00101010000000011111111111111111",
		"11111111111111000000000000000000",
		"00100100100111111111111111111111", -- 0x18F(399)  3. VLIW 
		"11111111111111111111111111111111",
		"11111111111000111000100001000011",
		"11111111111111111111111111111111", -- 0x192(402)  4. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x195(405)  5. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x198(408)  6. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x19B(411)  7. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x19E(414)  8. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x1A1(417)  9. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x1A4(420)  10. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x1A7(423)  11. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x1AA(426)  12. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x1AD(429)  13. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		"11111111111111111111111111111111", -- 0x1B0(432)  14. VLIW 
		"11111111111111111111111111111111",
		"11111111111111000000000000000000",
		--________________________________
		--==  Domain12 Header Parsing: [ Type: 1 (VLIW), lastFlag: 0, Next: 435, Vertical Mask: "10", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 390, VLIW end: 435, ICN begin: 511, ICN end: 511 ]
		--================================
		--
		"11111111110101111010110110110010", -- 0x1B3(435)  Domain_13, Type: ICN, Vert.Mask:2 "10" Horiz.Mask:2 "10",  *** PE[0,0] *** d1 INVERT ICN
		"11111111011011011011010111111111",
		"11111111111111111111000001111111",
		--________________________________
		--==  Domain13 Header Parsing: [ Type: 2 (ICN), lastFlag: 0, Next: 438, Vertical Mask: "10", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 511, VLIW end: 511, ICN begin: 437, ICN end: 438 ]
		--================================
		--
		"11111111110101111001111111111110", -- 0x1B6(438)  Domain_14, Type: ICN, LAST, Vert.Mask:1 "01" Horiz.Mask:2 "10",  *** PE[0,1] *** d2 INVERT ICN
		"11111111011100111011100011111111",
		"11111111111111111111111111000000",
		--________________________________
		--==  Domain14 Header Parsing: [ Type: 2 (ICN), lastFlag: 1, Next: 511, Vertical Mask: "01", Horizontal Mask: "10",
		--== VLIW Ratio: 3, ICN Ratio: 5, CountDown: 0, VLIW begin: 511, VLIW end: 511, ICN begin: 440, ICN end: 441 ]
		--================================
		--
		"11111111111111111111111111111111", -- 0x1B9(441)  Begin 71 Rest Memory Block(s)
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111",
		"11111111111111111111111111111111" -- 0x1FF(511)  End 71 Rest Memory Block(s)
	);

begin
	FPGA_SYN_CONFIG_MEM : IF FPGA_SYN GENERATE
		xilinx_data : process(clk, addr, we, d_in, ram) --, rst)	--== uncomment 1 of 4 for ASIC:


		begin
			if clk'event and clk = '1' then
				if we = '1' then        -- write enable

					ram(conv_integer(addr(ADDR_WIDTH - 1 downto 0))) <= d_in;

				else
					d_out <= ram(conv_integer(addr(ADDR_WIDTH - 1 downto 0)));

				end if;

			end if;

		end process xilinx_data;
	END GENERATE FPGA_SYN_CONFIG_MEM;

end Behavioral;
